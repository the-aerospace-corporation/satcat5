--------------------------------------------------------------------------
-- Copyright 2020-2024 The Aerospace Corporation.
-- This file is a part of SatCat5, licensed under CERN-OHL-W v2 or later.
--------------------------------------------------------------------------
--
-- SGMII port using the Xilinx Ethernet SGMII-PCS core
--
-- This module is a thin wrapper for a Xilinx SGMII IP core, "1G/2.5G Ethernet
-- PCS/PMA or SGMII", that uses a GTX SERDES to implement an SGMII connection.
--
-- Documentation for this IP core is in Xilinx document PG047:
-- https://www.xilinx.com/support/documentation/ip_documentation/gig_ethernet_pcs_pma/v16_1/pg047-gig-eth-pcs-pma.pdf
--
-- This block depends on the IP-core, which can be added to the Vivado project
-- by running "generate_sgmii_gtx.tcl" in the Xilinx projects folder and then
-- calling the newly-defined function(s) with various parameters.
--
-- To instantiate a single port:
--  * From the SatCat5 "project/vivado" folder:
--      * Run `source generate_sgmii_gtx.tcl`
--      * Run `generate_sgmii_gtx X0Y0`
--  * Instantiate a single "port_sgmii_gtx" block with SHARED_EN = true.
--
-- To instantiate multiple ports in the same quad:
--  * From a TCL console in the SatCat5 "project/vivado" folder:
--      * Run `source generate_sgmii_gtx.tcl`
--      * For 7-series parts:
--          * Run `generate_sgmii_gtx X0Y0 sgmii_gtx2 1`
--          * Run `generate_sgmii_gtx X0Y0 sgmii_gtx3 0`
--      * For Ultrascale and above:
--          * Run `generate_sgmii_gtx X0Y0 sgmii_gtx0 1`
--          * Run `generate_sgmii_gtx X0Y0 sgmii_gtx1 0`
--  * Instantiate the first "port_sgmii_gtx" block with SHARED_EN = true.
--  * Instantiate remaining "port_sgmii_gtx" block(s) with SHARED_EN = false.
--    Link each "shared_in" port to "shared_out" port on the first instance.
--  * For 7-series parts, also set SHARED_QPLL = true for all of the above.
--
-- For an SGMII port using regular GPIO, see "port_sgmii_gpio".
--

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;
use     work.common_functions.all;
use     work.common_primitives.all;
use     work.eth_frame_common.all;
use     work.ptp_types.all;
use     work.switch_types.all;

entity port_sgmii_gtx is
    generic (
    AUTONEG_EN  : boolean;          -- Enable or disable autonegotiation
    SHARED_EN   : boolean := true;  -- Does the IP-core include shared logic?
    SHARED_QPLL : boolean := false; -- Workaround for shared QPLL signals?
    VCONFIG     : vernier_config := VERNIER_DISABLED);
    port (
    -- External SGMII interfaces (direct to GTX pins)
    sgmii_rxp   : in  std_logic;
    sgmii_rxn   : in  std_logic;
    sgmii_txp   : out std_logic;
    sgmii_txn   : out std_logic;

    -- Generic internal port interfaces.
    prx_data    : out port_rx_m2s;
    ptx_data    : in  port_tx_s2m;
    ptx_ctrl    : out port_tx_m2s;
    port_shdn   : in  std_logic;

    -- Global reference for PTP timestamps, if enabled.
    ref_time    : in  port_timeref := PORT_TIMEREF_NULL;

    -- Shared-logic enabled?
    -- Note: 7-Series RefClk = 125 MHz, Ultrascale = Required RefClk frequency
    gtrefclk_p  : in  std_logic := '0'; -- GTX RefClk, 125MHz on 7 series
    gtrefclk_n  : in  std_logic := '0'; -- (Differential)
    shared_out  : out std_logic_vector(15 downto 0);

    -- Shared-logic disabled?
    shared_in   : in  std_logic_vector(15 downto 0) := (others => '0');

    -- Additional clocks.
    clkin_bufg  : in  std_logic;    -- IDELAYCTRL or DRP clock
    clkout_125  : out std_logic);   -- Optional 125 MHz output
end port_sgmii_gtx;

architecture port_sgmii_gtx of port_sgmii_gtx is

-- Component declaration for different variations on the black-box IP core.
-- Note: If shared-logic is enabled, then the "gtx0" variant is compatible
--   with all supported platforms. i.e., All undefined signals are outputs.
component sgmii_gtx0 is     -- Shared logic, no QPLL
    port(
    gtrefclk_p              : in  std_logic;
    gtrefclk_n              : in  std_logic;
    gtrefclk_out            : out std_logic;
    txp                     : out std_logic;
    txn                     : out std_logic;
    rxp                     : in std_logic;
    rxn                     : in std_logic;
    resetdone               : out std_logic;
    userclk_out             : out std_logic;
    userclk2_out            : out std_logic;
    rxuserclk_out           : out std_logic;
    rxuserclk2_out          : out std_logic;
    pma_reset_out           : out std_logic;
    mmcm_locked_out         : out std_logic;
    independent_clock_bufg  : in std_logic;
    sgmii_clk_r             : out std_logic;
    sgmii_clk_f             : out std_logic;
    sgmii_clk_en            : out std_logic;
    gmii_txd                : in std_logic_vector(7 downto 0);
    gmii_tx_en              : in std_logic;
    gmii_tx_er              : in std_logic;
    gmii_rxd                : out std_logic_vector(7 downto 0);
    gmii_rx_dv              : out std_logic;
    gmii_rx_er              : out std_logic;
    gmii_isolate            : out std_logic;
    configuration_vector    : in std_logic_vector(4 downto 0);
    speed_is_10_100         : in std_logic;
    speed_is_100            : in std_logic;
    status_vector           : out std_logic_vector(15 downto 0);
    reset                   : in std_logic;
    gtpowergood             : out std_logic;
    signal_detect           : in std_logic);
end component;

component sgmii_gtx1 is     -- No shared logic, no QPLL
    port(
    gtrefclk                : in std_logic;
    txp                     : out std_logic;
    txn                     : out std_logic;
    rxp                     : in std_logic;
    rxn                     : in std_logic;
    resetdone               : out std_logic;
    userclk                 : in std_logic;
    userclk2                : in std_logic;
    rxuserclk               : in std_logic;
    rxuserclk2              : in std_logic;
    pma_reset               : in std_logic;
    mmcm_locked             : in std_logic;
    independent_clock_bufg  : in std_logic;
    sgmii_clk_r             : out std_logic;
    sgmii_clk_f             : out std_logic;
    sgmii_clk_en            : out std_logic;
    gmii_txd                : in std_logic_vector(7 downto 0);
    gmii_tx_en              : in std_logic;
    gmii_tx_er              : in std_logic;
    gmii_rxd                : out std_logic_vector(7 downto 0);
    gmii_rx_dv              : out std_logic;
    gmii_rx_er              : out std_logic;
    gmii_isolate            : out std_logic;
    configuration_vector    : in std_logic_vector(4 downto 0);
    status_vector           : out std_logic_vector(15 downto 0);
    reset                   : in std_logic;
    signal_detect           : in std_logic);
end component;

component sgmii_gtx2 is     -- Shared logic, with QPLL
    port(
    gtrefclk_p              : in  std_logic;
    gtrefclk_n              : in  std_logic;
    gtrefclk_out            : out std_logic;
    gtrefclk_bufg_out       : out std_logic;
    txp                     : out std_logic;
    txn                     : out std_logic;
    rxp                     : in std_logic;
    rxn                     : in std_logic;
    resetdone               : out std_logic;
    userclk_out             : out std_logic;
    userclk2_out            : out std_logic;
    rxuserclk_out           : out std_logic;
    rxuserclk2_out          : out std_logic;
    pma_reset_out           : out std_logic;
    mmcm_locked_out         : out std_logic;
    independent_clock_bufg  : in std_logic;
    sgmii_clk_r             : out std_logic;
    sgmii_clk_f             : out std_logic;
    sgmii_clk_en            : out std_logic;
    gmii_txd                : in std_logic_vector(7 downto 0);
    gmii_tx_en              : in std_logic;
    gmii_tx_er              : in std_logic;
    gmii_rxd                : out std_logic_vector(7 downto 0);
    gmii_rx_dv              : out std_logic;
    gmii_rx_er              : out std_logic;
    gmii_isolate            : out std_logic;
    configuration_vector    : in std_logic_vector(4 downto 0);
    speed_is_10_100         : in std_logic;
    speed_is_100            : in std_logic;
    status_vector           : out std_logic_vector(15 downto 0);
    reset                   : in std_logic;
    signal_detect           : in std_logic;
    gt0_qplloutclk_out      : out std_logic;
    gt0_qplloutrefclk_out   : out std_logic);
end component;

component sgmii_gtx3 is     -- No shared logic, with QPLL
    port(
    gtrefclk                : in std_logic;
    gtrefclk_bufg           : in std_logic;
    txp                     : out std_logic;
    txn                     : out std_logic;
    rxp                     : in std_logic;
    rxn                     : in std_logic;
    resetdone               : out std_logic;
    userclk                 : in std_logic;
    userclk2                : in std_logic;
    rxuserclk               : in std_logic;
    rxuserclk2              : in std_logic;
    pma_reset               : in std_logic;
    mmcm_locked             : in std_logic;
    independent_clock_bufg  : in std_logic;
    sgmii_clk_r             : out std_logic;
    sgmii_clk_f             : out std_logic;
    sgmii_clk_en            : out std_logic;
    gmii_txd                : in std_logic_vector(7 downto 0);
    gmii_tx_en              : in std_logic;
    gmii_tx_er              : in std_logic;
    gmii_rxd                : out std_logic_vector(7 downto 0);
    gmii_rx_dv              : out std_logic;
    gmii_rx_er              : out std_logic;
    gmii_isolate            : out std_logic;
    configuration_vector    : in std_logic_vector(4 downto 0);
    status_vector           : out std_logic_vector(15 downto 0);
    reset                   : in std_logic;
    signal_detect           : in std_logic;
    gt0_qplloutclk_in       : in std_logic;
    gt0_qplloutrefclk_in    : in std_logic);
end component;

-- Control signals
signal txrx_pwren       : std_logic;
signal tx_pkten         : std_logic;
signal config_vec       : std_logic_vector(4 downto 0);
signal status_vec       : std_logic_vector(15 downto 0);
signal status_linkok    : std_logic;
signal status_sync      : std_logic;
signal status_disperr   : std_logic;
signal status_badsymb   : std_logic;
signal status_phyok     : std_logic;
signal aux_err_async    : std_logic;
signal aux_err_sync     : std_logic;

-- Receiver timestamp logic, if enabled.
signal txrx_reset       : std_logic := '0';
signal rx_treset        : std_logic := '0';
signal rx_tstamp        : tstamp_t := TSTAMP_DISABLED;
signal rx_tfreq         : tfreq_t := TFREQ_DISABLED;
signal rx_tvalid        : std_logic := '0';
signal tx_treset        : std_logic := '0';
signal tx_tstamp        : tstamp_t := TSTAMP_DISABLED;
signal tx_tfreq         : tfreq_t := TFREQ_DISABLED;
signal tx_tvalid        : std_logic := '0';

-- IP-core provides a quasi-GMII interface.
signal gmii_tx_clk      : std_logic;
signal gmii_tx_data     : byte_t;
signal gmii_tx_en       : std_logic;
signal gmii_tx_er       : std_logic;
signal gmii_rx_clk      : std_logic;
signal gmii_rx_data     : byte_t;
signal gmii_rx_dv       : std_logic;
signal gmii_rx_er       : std_logic;
signal gmii_status      : port_status_t;

-- Other signals relating to shared-logic crosslinking.
signal xil_gtrefclk     : std_logic;
signal xil_gtrefbuf     : std_logic;
signal xil_userclk      : std_logic;
signal xil_userclk2     : std_logic;
signal xil_rxuserclk    : std_logic;
signal xil_rxuserclk2   : std_logic;
signal xil_mmcm_locked  : std_logic;
signal xil_pma_reset    : std_logic;
signal xil_qpll_clk     : std_logic;
signal xil_qpll_ref     : std_logic;

begin

-- Add preambles to the outgoing data:
u_amble_tx : entity work.eth_preamble_tx
    port map(
    out_data    => gmii_tx_data,
    out_dv      => gmii_tx_en,
    out_err     => gmii_tx_er,
    tx_clk      => gmii_tx_clk,
    tx_pwren    => txrx_pwren,
    tx_pkten    => tx_pkten,
    tx_tstamp   => tx_tstamp,
    tx_tfreq    => tx_tfreq,
    tx_data     => ptx_data,
    tx_ctrl     => ptx_ctrl);

-- Receiver timestamp logic, if enabled.
-- TODO: This logic doesn't have visibility into the Xilinx SGMII IP core.
--  As a result, various internal delays will result in uncontrolled error.
--  The error will likely be an integer multiple of the bit period and may
--  be quasi-static on each reset.  The end-to-end result could be up to
--  +/- 100 nsec of uncorrectable bias.  Later versions should integrate
--  the core's PTP timestamps to correct this deficiency.
gen_tstamp : if VCONFIG.input_hz > 0 generate
    txrx_reset <= not xil_mmcm_locked;

    u_rx_treset : sync_reset
        port map(
        in_reset_p  => txrx_reset,
        out_reset_p => rx_treset,
        out_clk     => gmii_rx_clk);

    u_tx_treset : sync_reset
        port map(
        in_reset_p  => txrx_reset,
        out_reset_p => tx_treset,
        out_clk     => gmii_tx_clk);

    u_rx_tstamp : entity work.ptp_counter_sync
        generic map(
        VCONFIG     => VCONFIG,
        USER_CLK_HZ => 125_000_000)
        port map(
        ref_time    => ref_time,
        user_clk    => gmii_rx_clk,
        user_ctr    => rx_tstamp,
        user_freq   => rx_tfreq,
        user_lock   => rx_tvalid,
        user_rst_p  => rx_treset);

    u_tx_tstamp : entity work.ptp_counter_sync
        generic map(
        VCONFIG     => VCONFIG,
        USER_CLK_HZ => 125_000_000)
        port map(
        ref_time    => ref_time,
        user_clk    => gmii_tx_clk,
        user_ctr    => tx_tstamp,
        user_freq   => tx_tfreq,
        user_lock   => tx_tvalid,
        user_rst_p  => tx_treset);
end generate;

-- Remove preambles from the incoming data:
u_amble_rx : entity work.eth_preamble_rx
    port map(
    raw_clk     => gmii_rx_clk,
    raw_lock    => xil_mmcm_locked,
    raw_data    => gmii_rx_data,
    raw_dv      => gmii_rx_dv,
    raw_err     => gmii_rx_er,
    rate_word   => get_rate_word(1000),
    rx_tstamp   => rx_tstamp,
    rx_tfreq    => rx_tfreq,
    aux_err     => aux_err_sync,
    status      => gmii_status,
    rx_data     => prx_data);

-- Flush received data if we get an 8b/10b decode error.
aux_err_async <= xil_mmcm_locked and (status_disperr or status_badsymb);

u_errsync : sync_toggle2pulse
    generic map(RISING_ONLY => true)
    port map(
    in_toggle   => aux_err_async,
    out_strobe  => aux_err_sync,
    out_clk     => gmii_rx_clk);

-- Other control signals:
txrx_pwren  <= not port_shdn;
tx_pkten    <= xil_mmcm_locked and status_linkok;

config_vec <= (
    4 => bool2bit(AUTONEG_EN),  -- Enable/disable auto-negotation
    3 => '0',                   -- Normal GMII operation
    2 => port_shdn,             -- Power-down strobe
    1 => '0',                   -- Disable loopback
    0 => '0');                  -- Bidirectional mode

status_linkok   <= status_vec(0);   -- SGMII link ready for use
status_sync     <= status_vec(1);   -- 8b/10b initial sync
status_disperr  <= status_vec(5);   -- 8b/10b disparity error
status_badsymb  <= status_vec(6);   -- 8b/10b decode error
status_phyok    <= status_vec(7);   -- Attached PHY status, if applicable

gmii_status <= (
    0 => port_shdn,
    1 => xil_mmcm_locked,
    2 => status_sync,
    3 => status_linkok,
    4 => status_phyok,
    5 => rx_tvalid and tx_tvalid,
    others => '0');

-- Alias for specific clock signals:
clkout_125  <= xil_gtrefclk;
gmii_rx_clk <= xil_userclk2;
gmii_tx_clk <= xil_userclk2;

-- Drive or accept shared-logic signals.
-- Note: Using 10 of 16 bits; the rest are reserved for future expansion.
shared_out <= (
    0 => xil_gtrefclk,
    1 => xil_gtrefbuf,
    2 => xil_userclk,
    3 => xil_userclk2,
    4 => xil_rxuserclk,
    5 => xil_rxuserclk2,
    6 => xil_pma_reset,
    7 => xil_mmcm_locked,
    8 => xil_qpll_clk,
    9 => xil_qpll_ref,
    others => '0');

-- When SHARED_EN = True, gtrefclk, gtrefbuf, userclk, etc.
-- are output signals of sgmii_gtx IP core
-- when SHARED_EN = False, these signals are inputs
gen_shared : if not SHARED_EN generate
    xil_gtrefclk    <= shared_in(0);
    xil_gtrefbuf    <= shared_in(1);
    xil_userclk     <= shared_in(2);
    xil_userclk2    <= shared_in(3);
    xil_rxuserclk   <= shared_in(4);
    xil_rxuserclk2  <= shared_in(5);
    xil_pma_reset   <= shared_in(6);
    xil_mmcm_locked <= shared_in(7);
    xil_qpll_clk    <= shared_in(8);
    xil_qpll_ref    <= shared_in(9);
end generate;

-- Instantiate the selected variant of the IP-core.
gen_variant0 : if (SHARED_EN) and (not SHARED_QPLL) generate
    xil_gtrefbuf <= xil_gtrefclk;
    xil_qpll_clk <= '0';
    xil_qpll_ref <= '0';

    u_ipcore : sgmii_gtx0
        port map(
        gtrefclk_p              => gtrefclk_p,
        gtrefclk_n              => gtrefclk_n,
        gtrefclk_out            => xil_gtrefclk,    -- Internal 125 MHz
        txp                     => sgmii_txp,
        txn                     => sgmii_txn,
        rxp                     => sgmii_rxp,
        rxn                     => sgmii_rxn,
        resetdone               => open,
        userclk_out             => xil_userclk,     -- Tx 62.5 MHz
        userclk2_out            => xil_userclk2,    -- Tx 125 MHz
        rxuserclk_out           => xil_rxuserclk,   -- Rx 62.5 MHz
        rxuserclk2_out          => xil_rxuserclk2,  -- Rx 62.5 MHz
        pma_reset_out           => xil_pma_reset,
        mmcm_locked_out         => xil_mmcm_locked,
        independent_clock_bufg  => clkin_bufg,      -- Clock for control logic
        sgmii_clk_r             => open,            -- Line-rate Tx clock
        sgmii_clk_f             => open,
        sgmii_clk_en            => open,
        gmii_txd                => gmii_tx_data,    -- GMII Tx
        gmii_tx_en              => gmii_tx_en,
        gmii_tx_er              => gmii_tx_er,
        gmii_rxd                => gmii_rx_data,    -- GMII Rx
        gmii_rx_dv              => gmii_rx_dv,
        gmii_rx_er              => gmii_rx_er,
        gmii_isolate            => open,
        configuration_vector    => config_vec,      -- See PG047, Table 2-39
        speed_is_10_100         => '0',             -- Always 1000 Mbps
        speed_is_100            => '0',             -- Always 1000 Mbps
        status_vector           => status_vec,      -- See PG047, Table 2-41
        reset                   => port_shdn,       -- Reset the entire core
        gtpowergood             => open,
        signal_detect           => '1');
end generate;

gen_variant1 : if (not SHARED_EN) and (not SHARED_QPLL) generate
    u_ipcore : sgmii_gtx1
        port map(
        gtrefclk                => xil_gtrefclk,    -- Internal 125 MHz
        txp                     => sgmii_txp,
        txn                     => sgmii_txn,
        rxp                     => sgmii_rxp,
        rxn                     => sgmii_rxn,
        resetdone               => open,
        userclk                 => xil_userclk,     -- Tx 62.5 MHz
        userclk2                => xil_userclk2,    -- Tx 125 MHz
        rxuserclk               => xil_rxuserclk,   -- Rx 62.5 MHz
        rxuserclk2              => xil_rxuserclk2,  -- Rx 62.5 MHz
        pma_reset               => xil_pma_reset,
        mmcm_locked             => xil_mmcm_locked,
        independent_clock_bufg  => clkin_bufg,      -- Clock for control logic
        sgmii_clk_r             => open,            -- Line-rate Tx clock
        sgmii_clk_f             => open,
        sgmii_clk_en            => open,
        gmii_txd                => gmii_tx_data,    -- GMII Tx
        gmii_tx_en              => gmii_tx_en,
        gmii_tx_er              => gmii_tx_er,
        gmii_rxd                => gmii_rx_data,    -- GMII Rx
        gmii_rx_dv              => gmii_rx_dv,
        gmii_rx_er              => gmii_rx_er,
        gmii_isolate            => open,
        configuration_vector    => config_vec,      -- See PG047, Table 2-39
        status_vector           => status_vec,      -- See PG047, Table 2-41
        reset                   => port_shdn,       -- Reset the entire core
        signal_detect           => '1');
end generate;

gen_variant2 : if (SHARED_EN) and (SHARED_QPLL) generate
    u_ipcore : sgmii_gtx2
        port map(
        gtrefclk_p              => gtrefclk_p,
        gtrefclk_n              => gtrefclk_n,
        gtrefclk_out            => xil_gtrefclk,    -- Internal 125 MHz
        gtrefclk_bufg_out       => xil_gtrefbuf,
        txp                     => sgmii_txp,
        txn                     => sgmii_txn,
        rxp                     => sgmii_rxp,
        rxn                     => sgmii_rxn,
        resetdone               => open,
        userclk_out             => xil_userclk,     -- Tx 62.5 MHz
        userclk2_out            => xil_userclk2,    -- Tx 125 MHz
        rxuserclk_out           => xil_rxuserclk,   -- Rx 62.5 MHz
        rxuserclk2_out          => xil_rxuserclk2,  -- Rx 62.5 MHz
        pma_reset_out           => xil_pma_reset,
        mmcm_locked_out         => xil_mmcm_locked,
        independent_clock_bufg  => clkin_bufg,      -- Clock for control logic
        sgmii_clk_r             => open,            -- Line-rate Tx clock
        sgmii_clk_f             => open,
        sgmii_clk_en            => open,
        gmii_txd                => gmii_tx_data,    -- GMII Tx
        gmii_tx_en              => gmii_tx_en,
        gmii_tx_er              => gmii_tx_er,
        gmii_rxd                => gmii_rx_data,    -- GMII Rx
        gmii_rx_dv              => gmii_rx_dv,
        gmii_rx_er              => gmii_rx_er,
        gmii_isolate            => open,
        configuration_vector    => config_vec,      -- See PG047, Table 2-39
        speed_is_10_100         => '0',             -- Always 1000 Mbps
        speed_is_100            => '0',             -- Always 1000 Mbps
        status_vector           => status_vec,      -- See PG047, Table 2-41
        reset                   => port_shdn,       -- Reset the entire core
        signal_detect           => '1',
        gt0_qplloutclk_out      => xil_qpll_clk,
        gt0_qplloutrefclk_out   => xil_qpll_ref);
end generate;

gen_variant3 : if (not SHARED_EN) and (SHARED_QPLL) generate
    u_ipcore : sgmii_gtx3
        port map(
        gtrefclk                => xil_gtrefclk,    -- Internal 125 MHz
        gtrefclk_bufg           => xil_gtrefbuf,
        txp                     => sgmii_txp,
        txn                     => sgmii_txn,
        rxp                     => sgmii_rxp,
        rxn                     => sgmii_rxn,
        resetdone               => open,
        userclk                 => xil_userclk,     -- Tx 62.5 MHz
        userclk2                => xil_userclk2,    -- Tx 125 MHz
        rxuserclk               => xil_rxuserclk,   -- Rx 62.5 MHz
        rxuserclk2              => xil_rxuserclk2,  -- Rx 62.5 MHz
        pma_reset               => xil_pma_reset,
        mmcm_locked             => xil_mmcm_locked,
        independent_clock_bufg  => clkin_bufg,      -- Clock for control logic
        sgmii_clk_r             => open,            -- Line-rate Tx clock
        sgmii_clk_f             => open,
        sgmii_clk_en            => open,
        gmii_txd                => gmii_tx_data,    -- GMII Tx
        gmii_tx_en              => gmii_tx_en,
        gmii_tx_er              => gmii_tx_er,
        gmii_rxd                => gmii_rx_data,    -- GMII Rx
        gmii_rx_dv              => gmii_rx_dv,
        gmii_rx_er              => gmii_rx_er,
        gmii_isolate            => open,
        configuration_vector    => config_vec,      -- See PG047, Table 2-39
        status_vector           => status_vec,      -- See PG047, Table 2-41
        reset                   => port_shdn,       -- Reset the entire core
        signal_detect           => '1',
        gt0_qplloutclk_in       => xil_qpll_clk,
        gt0_qplloutrefclk_in    => xil_qpll_ref);
end generate;

end port_sgmii_gtx;
