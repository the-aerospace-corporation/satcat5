--------------------------------------------------------------------------
-- Copyright 2025 The Aerospace Corporation.
-- This file is a part of SatCat5, licensed under CERN-OHL-W v2 or later.
--------------------------------------------------------------------------
-- Microsemi SGMII port using a standard I/O pin via IOD-CDR primitives.
--
-- UNTESTED as of March 2025 due to issues with the PolarFire Eval Kit PHY.
--
-- Requires Mircosemi IP generated by project/libero/ipcores/sgmii_gpio.tcl.
--
-- This module uses the PF_IOD_CDR and PF_IOD_CDR_CCC IP cores which handle CDR
-- and phase/voltage/temp compensation for the RX line using features built into
-- digital I/O (IOD) pins of the FPGA. This core adds required encode/decode and
-- adapts the interface to act as one or more ports on a SatCat5 switch. Any
-- number of lanes can be generated - all will share a single set of generated
-- clocks from PF_IOD_CDR_CCC as recommended by Microsemi.
--
-- See also Microsemi documentation:
--  * AN4623: 1G Ethernet Using Transceiver
--  * UG0687: 1G Ethernet Solutions User Guide
--

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;
use     work.common_primitives.all;
use     work.ptp_types.all;
use     work.switch_types.all;

entity port_sgmii_gpio is
generic (
    LANES       : integer := 1;         -- Number of port lanes to generate
    SHAKE_WAIT  : boolean := false;     -- Wait for MAC/PHY handshake?
    VCONFIG     : vernier_config := VERNIER_DISABLED);
port (
    -- External SGMII interfaces (direct to FPGA pins)
    sgmii_rxp   : in  std_logic_vector(LANES-1 downto 0);
    sgmii_rxn   : in  std_logic_vector(LANES-1 downto 0);
    sgmii_txp   : out std_logic_vector(LANES-1 downto 0);
    sgmii_txn   : out std_logic_vector(LANES-1 downto 0);

    -- Global reference for PTP timestamps, if enabled.
    -- TODO: This block currently does not support PTP, this is left as a stub.
    ref_time    : in  port_timeref := PORT_TIMEREF_NULL;

    -- Generic internal port interfaces.
    prx_data    : out array_rx_m2s(LANES-1 downto 0);
    ptx_data    : in  array_tx_s2m(LANES-1 downto 0);
    ptx_ctrl    : out array_tx_m2s(LANES-1 downto 0);
    port_shdn   : in  std_logic_vector(LANES-1 downto 0);
    port_test   : in  std_logic_vector(LANES-1 downto 0) := (others => '0');

    -- Reference clocks and reset.
    clk_125     : in  std_logic;
    stream_start: in  std_logic;
    reset_p     : in  std_logic);
end port_sgmii_gpio;

architecture microsemi of port_sgmii_gpio is

-- Clocking and reset.
signal reset_n          : std_logic;
signal tx_clk           : std_logic;
signal rx_clk           : std_logic_vector(LANES-1 downto 0);

-- IOD_CDR clocking signals, routed from clocking to all instances.
signal cdr_start        : std_logic;
signal dll_delay_code   : std_logic_vector(6 downto 0);
signal dll_lock         : std_logic;
signal dll_valid_code   : std_logic;
signal hs_io_clk_0      : std_logic;
signal hs_io_clk_90     : std_logic;
signal hs_io_clk_180    : std_logic;
signal hs_io_clk_270    : std_logic;
signal hs_io_clk_pause  : std_logic;
signal pll_lock         : std_logic;
signal tx_clk_to_cdr    : std_logic; -- Route to IOD_CDR IP, tx_clk for logic.

-- TX/RX parallel data signals.
signal tx_data10        : std_logic_vector(10*LANES-1 downto 0);
signal rx_data10        : std_logic_vector(10*LANES-1 downto 0);
signal rx_valid         : std_logic_vector(LANES-1 downto 0);

-- Microsemi IP: PF_IOD_CDR_CCC:2.1.111
component PF_IOD_CDR_CCC_SGMII
port (
    ARST_N          : in  std_logic;
    REF_CLK         : in  std_logic;
    CDR_START       : out std_logic;
    DLL_DELAY_CODE  : out std_logic_vector(6 downto 0);
    DLL_LOCK        : out std_logic;
    DLL_VALID_CODE  : out std_logic;
    HS_IO_CLK_0     : out std_logic;
    HS_IO_CLK_90    : out std_logic;
    HS_IO_CLK_180   : out std_logic;
    HS_IO_CLK_270   : out std_logic;
    HS_IO_CLK_PAUSE : out std_logic;
    PLL_LOCK        : out std_logic;
    TX_CLK_G        : out std_logic;
    TX_CLK_G_TO_CDR : out std_logic);
end component;

-- Microsemi IP: PF_IOD_CDR:2.4.105
component PF_IOD_CDR_SGMII
port (
    CDR_START       : in  std_logic;
    DLL_DELAY_CODE  : in  std_logic_vector(6 downto 0);
    DLL_LOCK        : in  std_logic;
    DLL_VALID_CODE  : in  std_logic;
    HS_IO_CLK_0     : in  std_logic;
    HS_IO_CLK_90    : in  std_logic;
    HS_IO_CLK_180   : in  std_logic;
    HS_IO_CLK_270   : in  std_logic;
    HS_IO_CLK_PAUSE : in  std_logic;
    PLL_LOCK        : in  std_logic;
    RST_N           : in  std_logic;
    RX_N            : in  std_logic;
    RX_P            : in  std_logic;
    STREAM_START    : in  std_logic;
    TX_CLK_G        : in  std_logic;
    TX_DATA         : in  std_logic_vector(9 downto 0);
    RX_CLK_R        : out std_logic;
    RX_DATA         : out std_logic_vector(9 downto 0);
    RX_VAL          : out std_logic;
    TX_N            : out std_logic;
    TX_P            : out std_logic);
end component;

begin

-- Clocking and reset.
reset_n <= not reset_p;

-- Common clocking infrastructure for all cores.
u_iod_cdr_ccc : PF_IOD_CDR_CCC_SGMII
port map (
    ARST_N          => reset_n,
    REF_CLK         => clk_125,
    CDR_START       => cdr_start,
    DLL_DELAY_CODE  => dll_delay_code,
    DLL_LOCK        => dll_lock,
    DLL_VALID_CODE  => dll_valid_code,
    HS_IO_CLK_0     => hs_io_clk_0,
    HS_IO_CLK_90    => hs_io_clk_90,
    HS_IO_CLK_180   => hs_io_clk_180,
    HS_IO_CLK_270   => hs_io_clk_270,
    HS_IO_CLK_PAUSE => hs_io_clk_pause,
    PLL_LOCK        => pll_lock,
    TX_CLK_G        => tx_clk,
    TX_CLK_G_TO_CDR => tx_clk_to_cdr);

-- Generate one or more IOD_CDR instances and route to port_smgii_common.
gen_lanes : for n in 0 to LANES-1 generate

    -- Performs clock and data recovery, outputs ten-bit interface (TBI).
    -- Note: UG0686 very specifically calls out that STREAM_START must be
    -- controlled to go high to indicate the incoming data stream is valid and
    -- may NOT be tied high. Use port_sgmii_common's decoder lock for this
    -- validation. AN4623 sets up a small state machine to look for transitions
    -- in RX_DATA, so this is probably fine.
    u_iod_cdr : PF_IOD_CDR_SGMII
    port map (
        CDR_START       => cdr_start,
        DLL_DELAY_CODE  => dll_delay_code,
        DLL_LOCK        => dll_lock,
        DLL_VALID_CODE  => dll_valid_code,
        HS_IO_CLK_0     => hs_io_clk_0,
        HS_IO_CLK_90    => hs_io_clk_90,
        HS_IO_CLK_180   => hs_io_clk_180,
        HS_IO_CLK_270   => hs_io_clk_270,
        HS_IO_CLK_PAUSE => hs_io_clk_pause,
        PLL_LOCK        => pll_lock,
        RST_N           => reset_n,
        RX_N            => sgmii_rxn(n),
        RX_P            => sgmii_rxp(n),
        STREAM_START    => stream_start,
        TX_CLK_G        => tx_clk_to_cdr,
        TX_DATA         => tx_data10((n+1)*10-1 downto n*10),
        RX_CLK_R        => rx_clk(n),
        RX_DATA         => rx_data10((n+1)*10-1 downto n*10),
        RX_VAL          => rx_valid(n),
        TX_N            => sgmii_txn(n),
        TX_P            => sgmii_txp(n));

    -- Handles SGMII logic including 8b/10b, handshaking, and preambles.
    -- TODO: All timestamping (rx/tx_tstamp/tfreq/tvalid) will need to be routed
    -- to PTP blocks (ptp_counter_sync) once this core is up.
    u_if : entity work.port_sgmii_common
    generic map (
        SHAKE_WAIT  => SHAKE_WAIT)
    port map (
        tx_clk      => tx_clk,
        tx_cken     => pll_lock,
        tx_data     => tx_data10((n+1)*10-1 downto n*10),
        tx_tstamp   => TSTAMP_DISABLED,
        tx_tfreq    => TFREQ_DISABLED,
        tx_tvalid   => '0',
        port_test   => port_test(n),
        rx_clk      => rx_clk(n),
        rx_cken     => pll_lock,
        rx_lock     => rx_valid(n),
        rx_data     => rx_data10((n+1)*10-1 downto n*10),
        rx_tstamp   => TSTAMP_DISABLED,
        rx_tfreq    => TFREQ_DISABLED,
        rx_tvalid   => '0',
        prx_data    => prx_data(n),
        ptx_data    => ptx_data(n),
        ptx_ctrl    => ptx_ctrl(n),
        reset_p     => reset_p);
end generate;

end microsemi;
