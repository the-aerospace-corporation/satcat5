--------------------------------------------------------------------------
-- Copyright 2019 The Aerospace Corporation
--
-- This file is part of SatCat5.
--
-- SatCat5 is free software: you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License as published by the
-- Free Software Foundation, either version 3 of the License, or (at your
-- option) any later version.
--
-- SatCat5 is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU Lesser General Public
-- License for more details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with SatCat5.  If not, see <https://www.gnu.org/licenses/>.
--------------------------------------------------------------------------
--
-- Constants for the Ethernet 8b/10b encoder
--
-- This package defines a large lookup table for the 8b/10b encoder.
-- It is separated from the main file, eth_enc8b10b, for better readability.
--
-- The index to the table is the combined code state:
--   * Bit 9: Is this a control token ('1') or a data token ('0')?
--   * Bit 8: Is the running disparity positive ('1') or negative ('0')?
--   * Bit 7-0: The octet value to be encoded ("H" in MSB).
--
-- The result is as follows:
--   * Bit 10: Set if the running disparity should be toggled.
--   * Bits 9-0: The output token ("abcdefghij", "a" in MSB).
--
-- The resulting 1024x11 ROM fits inside an 18 kbit BRAM.  Since it is read-only,
-- and each BRAM has two read ports, two 8b/10b encoders may share a single BRAM.
--
-- The table contents are generated by the MATLAB script "make_8b10b_table.m".
--
-- For more information, refer to:
--   IEEE 802.3 Section 3.36, Table 36-1 and 36-2.
--   http://standards.ieee.org/getieee802/802.3.html
--   https://ieeexplore.ieee.org/xpl/mostRecentIssue.jsp?punumber=7428774
--

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

package eth_enc8b10b_table is
    subtype rom_index is integer range 0 to 1023;
    subtype rom_word is std_logic_vector(10 downto 0);
    type rom_array is array(0 to 1023) of rom_word;

    constant ENC_TABLE : rom_array := (
    "01001101010",
    "00111001010",
    "01011001010",
    "11100010111",
    "01101001010",
    "11010010111",
    "10110010111",
    "11110010101",
    "01110001010",
    "11001010111",
    "10101010111",
    "11101010101",
    "10011010111",
    "11011010101",
    "10111010101",
    "00101101010",
    "00110101010",
    "11000110111",
    "10100110111",
    "11100110101",
    "10010110111",
    "11010110101",
    "10110110101",
    "01110101000",
    "01100101010",
    "11001110101",
    "10101110101",
    "01101101000",
    "10011110101",
    "01011101000",
    "00111101000",
    "01010101010",
    "11001110011",
    "10111010011",
    "11011010011",
    "01100010011",
    "11101010011",
    "01010010011",
    "00110010011",
    "01110010001",
    "11110010011",
    "01001010011",
    "00101010011",
    "01101010001",
    "00011010011",
    "01011010001",
    "00111010001",
    "10101110011",
    "10110110011",
    "01000110011",
    "00100110011",
    "01100110001",
    "00010110011",
    "01010110001",
    "00110110001",
    "11110110001",
    "11100110011",
    "01001110001",
    "00101110001",
    "11101110001",
    "00011110001",
    "11011110001",
    "10111110001",
    "11010110011",
    "11001101011",
    "10111001011",
    "11011001011",
    "01100001011",
    "11101001011",
    "01010001011",
    "00110001011",
    "01110001001",
    "11110001011",
    "01001001011",
    "00101001011",
    "01101001001",
    "00011001011",
    "01011001001",
    "00111001001",
    "10101101011",
    "10110101011",
    "01000101011",
    "00100101011",
    "01100101001",
    "00010101011",
    "01010101001",
    "00110101001",
    "11110101001",
    "11100101011",
    "01001101001",
    "00101101001",
    "11101101001",
    "00011101001",
    "11011101001",
    "10111101001",
    "11010101011",
    "11001100111",
    "10111000111",
    "11011000111",
    "01100011010",
    "11101000111",
    "01010011010",
    "00110011010",
    "01110011000",
    "11110000111",
    "01001011010",
    "00101011010",
    "01101011000",
    "00011011010",
    "01011011000",
    "00111011000",
    "10101100111",
    "10110100111",
    "01000111010",
    "00100111010",
    "01100111000",
    "00010111010",
    "01010111000",
    "00110111000",
    "11110100101",
    "11100100111",
    "01001111000",
    "00101111000",
    "11101100101",
    "00011111000",
    "11011100101",
    "10111100101",
    "11010100111",
    "01001100110",
    "00111000110",
    "01011000110",
    "11100011011",
    "01101000110",
    "11010011011",
    "10110011011",
    "11110011001",
    "01110000110",
    "11001011011",
    "10101011011",
    "11101011001",
    "10011011011",
    "11011011001",
    "10111011001",
    "00101100110",
    "00110100110",
    "11000111011",
    "10100111011",
    "11100111001",
    "10010111011",
    "11010111001",
    "10110111001",
    "01110100100",
    "01100100110",
    "11001111001",
    "10101111001",
    "01101100100",
    "10011111001",
    "01011100100",
    "00111100100",
    "01010100110",
    "11001110110",
    "10111010110",
    "11011010110",
    "01100010110",
    "11101010110",
    "01010010110",
    "00110010110",
    "01110010100",
    "11110010110",
    "01001010110",
    "00101010110",
    "01101010100",
    "00011010110",
    "01011010100",
    "00111010100",
    "10101110110",
    "10110110110",
    "01000110110",
    "00100110110",
    "01100110100",
    "00010110110",
    "01010110100",
    "00110110100",
    "11110110100",
    "11100110110",
    "01001110100",
    "00101110100",
    "11101110100",
    "00011110100",
    "11011110100",
    "10111110100",
    "11010110110",
    "11001101110",
    "10111001110",
    "11011001110",
    "01100001110",
    "11101001110",
    "01010001110",
    "00110001110",
    "01110001100",
    "11110001110",
    "01001001110",
    "00101001110",
    "01101001100",
    "00011001110",
    "01011001100",
    "00111001100",
    "10101101110",
    "10110101110",
    "01000101110",
    "00100101110",
    "01100101100",
    "00010101110",
    "01010101100",
    "00110101100",
    "11110101100",
    "11100101110",
    "01001101100",
    "00101101100",
    "11101101100",
    "00011101100",
    "11011101100",
    "10111101100",
    "11010101110",
    "01001100011",
    "00111000011",
    "01011000011",
    "11100011110",
    "01101000011",
    "11010011110",
    "10110011110",
    "11110011100",
    "01110000011",
    "11001011110",
    "10101011110",
    "11101011100",
    "10011011110",
    "11011011100",
    "10111011100",
    "00101100011",
    "00110100011",
    "11000101111",
    "10100101111",
    "11100111100",
    "10010101111",
    "11010111100",
    "10110111100",
    "01110100001",
    "01100100011",
    "11001111100",
    "10101111100",
    "01101100001",
    "10011111100",
    "01011100001",
    "00111100001",
    "01010100011",
    "00110010101",
    "01000110101",
    "00100110101",
    "11100001010",
    "00010110101",
    "11010001010",
    "10110001010",
    "10001101010",
    "00001110101",
    "11001001010",
    "10101001010",
    "11101001000",
    "10011001010",
    "11011001000",
    "10111001000",
    "01010010101",
    "01001010101",
    "11000101010",
    "10100101010",
    "11100101000",
    "10010101010",
    "11010101000",
    "10110101000",
    "00001010111",
    "00011010101",
    "11001101000",
    "10101101000",
    "00010010111",
    "10011101000",
    "00100010111",
    "01000010111",
    "00101010101",
    "10110010001",
    "11000110001",
    "10100110001",
    "01100010011",
    "10010110001",
    "01010010011",
    "00110010011",
    "00001110011",
    "10001110001",
    "01001010011",
    "00101010011",
    "01101010001",
    "00011010011",
    "01011010001",
    "00111010001",
    "11010010001",
    "11001010001",
    "01000110011",
    "00100110011",
    "01100110001",
    "00010110011",
    "01010110001",
    "00110110001",
    "10001010011",
    "10011010001",
    "01001110001",
    "00101110001",
    "10010010011",
    "00011110001",
    "10100010011",
    "11000010011",
    "10101010001",
    "10110001001",
    "11000101001",
    "10100101001",
    "01100001011",
    "10010101001",
    "01010001011",
    "00110001011",
    "00001101011",
    "10001101001",
    "01001001011",
    "00101001011",
    "01101001001",
    "00011001011",
    "01011001001",
    "00111001001",
    "11010001001",
    "11001001001",
    "01000101011",
    "00100101011",
    "01100101001",
    "00010101011",
    "01010101001",
    "00110101001",
    "10001001011",
    "10011001001",
    "01001101001",
    "00101101001",
    "10010001011",
    "00011101001",
    "10100001011",
    "11000001011",
    "10101001001",
    "10110011000",
    "11000111000",
    "10100111000",
    "01100000111",
    "10010111000",
    "01010000111",
    "00110000111",
    "00001100111",
    "10001111000",
    "01001000111",
    "00101000111",
    "01101000101",
    "00011000111",
    "01011000101",
    "00111000101",
    "11010011000",
    "11001011000",
    "01000100111",
    "00100100111",
    "01100100101",
    "00010100111",
    "01010100101",
    "00110100101",
    "10001011010",
    "10011011000",
    "01001100101",
    "00101100101",
    "10010011010",
    "00011100101",
    "10100011010",
    "11000011010",
    "10101011000",
    "00110011001",
    "01000111001",
    "00100111001",
    "11100000110",
    "00010111001",
    "11010000110",
    "10110000110",
    "10001100110",
    "00001111001",
    "11001000110",
    "10101000110",
    "11101000100",
    "10011000110",
    "11011000100",
    "10111000100",
    "01010011001",
    "01001011001",
    "11000100110",
    "10100100110",
    "11100100100",
    "10010100110",
    "11010100100",
    "10110100100",
    "00001011011",
    "00011011001",
    "11001100100",
    "10101100100",
    "00010011011",
    "10011100100",
    "00100011011",
    "01000011011",
    "00101011001",
    "10110010100",
    "11000110100",
    "10100110100",
    "01100010110",
    "10010110100",
    "01010010110",
    "00110010110",
    "00001110110",
    "10001110100",
    "01001010110",
    "00101010110",
    "01101010100",
    "00011010110",
    "01011010100",
    "00111010100",
    "11010010100",
    "11001010100",
    "01000110110",
    "00100110110",
    "01100110100",
    "00010110110",
    "01010110100",
    "00110110100",
    "10001010110",
    "10011010100",
    "01001110100",
    "00101110100",
    "10010010110",
    "00011110100",
    "10100010110",
    "11000010110",
    "10101010100",
    "10110001100",
    "11000101100",
    "10100101100",
    "01100001110",
    "10010101100",
    "01010001110",
    "00110001110",
    "00001101110",
    "10001101100",
    "01001001110",
    "00101001110",
    "01101001100",
    "00011001110",
    "01011001100",
    "00111001100",
    "11010001100",
    "11001001100",
    "01000101110",
    "00100101110",
    "01100101100",
    "00010101110",
    "01010101100",
    "00110101100",
    "10001001110",
    "10011001100",
    "01001101100",
    "00101101100",
    "10010001110",
    "00011101100",
    "10100001110",
    "11000001110",
    "10101001100",
    "00110011100",
    "01000111100",
    "00100111100",
    "11100000011",
    "00010111100",
    "11010000011",
    "10110000011",
    "10001100011",
    "00001111100",
    "11001000011",
    "10101000011",
    "11101010000",
    "10011000011",
    "11011010000",
    "10111010000",
    "01010011100",
    "01001011100",
    "11000100011",
    "10100100011",
    "11100100001",
    "10010100011",
    "11010100001",
    "10110100001",
    "00001011110",
    "00011011100",
    "11001100001",
    "10101100001",
    "00010011110",
    "10011100001",
    "00100011110",
    "01000011110",
    "00101011100",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00011101010",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "10011110011",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "10011101011",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "10011100111",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00011100110",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "10011110110",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "10011101110",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "01110110000",
    "00111110000",
    "00111110000",
    "00111110000",
    "01101110000",
    "00011110010",
    "01011110000",
    "00111110000",
    "00111110000",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01100010101",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "11100001100",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "11100010100",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "11100011000",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01100011001",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "11100001001",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "11100010001",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "00001001111",
    "01000001111",
    "01000001111",
    "01000001111",
    "00010001111",
    "01100001101",
    "00100001111",
    "01000001111",
    "01000001111");
end package;
